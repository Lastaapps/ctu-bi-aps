`default_nettype none
module processor( input i_clk, _reset,
                  output [31:0] o_PC,
                  input  [31:0] i_instruction,
                  output o_WE,
                  output [31:0] o_address_to_mem,
                  output [31:0] o_data_to_mem,
                  input  [31:0] i_data_from_mem
                );


endmodule
`default_nettype wire
